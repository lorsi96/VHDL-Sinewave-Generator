library ieee;
use ieee.std_logic_1164.all;
use IEEE.numeric_std.all;

entity sine_lut is
    port(
        address_in: in std_logic_vector(9 downto 0);
        data_out: out std_logic_vector(7 downto 0)
    );
end sine_lut;

architecture sine_lut_arch of sine_lut is
begin
    process(address_in) is
        begin
            case address_in is
                when "0000000000" => data_out <= "01111111"; -- 0x7f
                when "0000000001" => data_out <= "10000000"; -- 0x80
                when "0000000010" => data_out <= "10000001"; -- 0x81
                when "0000000011" => data_out <= "10000010"; -- 0x82
                when "0000000100" => data_out <= "10000011"; -- 0x83
                when "0000000101" => data_out <= "10000011"; -- 0x83
                when "0000000110" => data_out <= "10000100"; -- 0x84
                when "0000000111" => data_out <= "10000101"; -- 0x85
                when "0000001000" => data_out <= "10000110"; -- 0x86
                when "0000001001" => data_out <= "10000111"; -- 0x87
                when "0000001010" => data_out <= "10000111"; -- 0x87
                when "0000001011" => data_out <= "10001000"; -- 0x88
                when "0000001100" => data_out <= "10001001"; -- 0x89
                when "0000001101" => data_out <= "10001010"; -- 0x8a
                when "0000001110" => data_out <= "10001010"; -- 0x8a
                when "0000001111" => data_out <= "10001011"; -- 0x8b
                when "0000010000" => data_out <= "10001100"; -- 0x8c
                when "0000010001" => data_out <= "10001101"; -- 0x8d
                when "0000010010" => data_out <= "10001110"; -- 0x8e
                when "0000010011" => data_out <= "10001110"; -- 0x8e
                when "0000010100" => data_out <= "10001111"; -- 0x8f
                when "0000010101" => data_out <= "10010000"; -- 0x90
                when "0000010110" => data_out <= "10010001"; -- 0x91
                when "0000010111" => data_out <= "10010010"; -- 0x92
                when "0000011000" => data_out <= "10010010"; -- 0x92
                when "0000011001" => data_out <= "10010011"; -- 0x93
                when "0000011010" => data_out <= "10010100"; -- 0x94
                when "0000011011" => data_out <= "10010101"; -- 0x95
                when "0000011100" => data_out <= "10010101"; -- 0x95
                when "0000011101" => data_out <= "10010110"; -- 0x96
                when "0000011110" => data_out <= "10010111"; -- 0x97
                when "0000011111" => data_out <= "10011000"; -- 0x98
                when "0000100000" => data_out <= "10011000"; -- 0x98
                when "0000100001" => data_out <= "10011001"; -- 0x99
                when "0000100010" => data_out <= "10011010"; -- 0x9a
                when "0000100011" => data_out <= "10011011"; -- 0x9b
                when "0000100100" => data_out <= "10011100"; -- 0x9c
                when "0000100101" => data_out <= "10011100"; -- 0x9c
                when "0000100110" => data_out <= "10011101"; -- 0x9d
                when "0000100111" => data_out <= "10011110"; -- 0x9e
                when "0000101000" => data_out <= "10011111"; -- 0x9f
                when "0000101001" => data_out <= "10011111"; -- 0x9f
                when "0000101010" => data_out <= "10100000"; -- 0xa0
                when "0000101011" => data_out <= "10100001"; -- 0xa1
                when "0000101100" => data_out <= "10100010"; -- 0xa2
                when "0000101101" => data_out <= "10100010"; -- 0xa2
                when "0000101110" => data_out <= "10100011"; -- 0xa3
                when "0000101111" => data_out <= "10100100"; -- 0xa4
                when "0000110000" => data_out <= "10100101"; -- 0xa5
                when "0000110001" => data_out <= "10100101"; -- 0xa5
                when "0000110010" => data_out <= "10100110"; -- 0xa6
                when "0000110011" => data_out <= "10100111"; -- 0xa7
                when "0000110100" => data_out <= "10101000"; -- 0xa8
                when "0000110101" => data_out <= "10101000"; -- 0xa8
                when "0000110110" => data_out <= "10101001"; -- 0xa9
                when "0000110111" => data_out <= "10101010"; -- 0xaa
                when "0000111000" => data_out <= "10101011"; -- 0xab
                when "0000111001" => data_out <= "10101011"; -- 0xab
                when "0000111010" => data_out <= "10101100"; -- 0xac
                when "0000111011" => data_out <= "10101101"; -- 0xad
                when "0000111100" => data_out <= "10101110"; -- 0xae
                when "0000111101" => data_out <= "10101110"; -- 0xae
                when "0000111110" => data_out <= "10101111"; -- 0xaf
                when "0000111111" => data_out <= "10110000"; -- 0xb0
                when "0001000000" => data_out <= "10110001"; -- 0xb1
                when "0001000001" => data_out <= "10110001"; -- 0xb1
                when "0001000010" => data_out <= "10110010"; -- 0xb2
                when "0001000011" => data_out <= "10110011"; -- 0xb3
                when "0001000100" => data_out <= "10110011"; -- 0xb3
                when "0001000101" => data_out <= "10110100"; -- 0xb4
                when "0001000110" => data_out <= "10110101"; -- 0xb5
                when "0001000111" => data_out <= "10110110"; -- 0xb6
                when "0001001000" => data_out <= "10110110"; -- 0xb6
                when "0001001001" => data_out <= "10110111"; -- 0xb7
                when "0001001010" => data_out <= "10111000"; -- 0xb8
                when "0001001011" => data_out <= "10111000"; -- 0xb8
                when "0001001100" => data_out <= "10111001"; -- 0xb9
                when "0001001101" => data_out <= "10111010"; -- 0xba
                when "0001001110" => data_out <= "10111011"; -- 0xbb
                when "0001001111" => data_out <= "10111011"; -- 0xbb
                when "0001010000" => data_out <= "10111100"; -- 0xbc
                when "0001010001" => data_out <= "10111101"; -- 0xbd
                when "0001010010" => data_out <= "10111101"; -- 0xbd
                when "0001010011" => data_out <= "10111110"; -- 0xbe
                when "0001010100" => data_out <= "10111111"; -- 0xbf
                when "0001010101" => data_out <= "10111111"; -- 0xbf
                when "0001010110" => data_out <= "11000000"; -- 0xc0
                when "0001010111" => data_out <= "11000001"; -- 0xc1
                when "0001011000" => data_out <= "11000001"; -- 0xc1
                when "0001011001" => data_out <= "11000010"; -- 0xc2
                when "0001011010" => data_out <= "11000011"; -- 0xc3
                when "0001011011" => data_out <= "11000011"; -- 0xc3
                when "0001011100" => data_out <= "11000100"; -- 0xc4
                when "0001011101" => data_out <= "11000101"; -- 0xc5
                when "0001011110" => data_out <= "11000101"; -- 0xc5
                when "0001011111" => data_out <= "11000110"; -- 0xc6
                when "0001100000" => data_out <= "11000111"; -- 0xc7
                when "0001100001" => data_out <= "11000111"; -- 0xc7
                when "0001100010" => data_out <= "11001000"; -- 0xc8
                when "0001100011" => data_out <= "11001001"; -- 0xc9
                when "0001100100" => data_out <= "11001001"; -- 0xc9
                when "0001100101" => data_out <= "11001010"; -- 0xca
                when "0001100110" => data_out <= "11001011"; -- 0xcb
                when "0001100111" => data_out <= "11001011"; -- 0xcb
                when "0001101000" => data_out <= "11001100"; -- 0xcc
                when "0001101001" => data_out <= "11001100"; -- 0xcc
                when "0001101010" => data_out <= "11001101"; -- 0xcd
                when "0001101011" => data_out <= "11001110"; -- 0xce
                when "0001101100" => data_out <= "11001110"; -- 0xce
                when "0001101101" => data_out <= "11001111"; -- 0xcf
                when "0001101110" => data_out <= "11010000"; -- 0xd0
                when "0001101111" => data_out <= "11010000"; -- 0xd0
                when "0001110000" => data_out <= "11010001"; -- 0xd1
                when "0001110001" => data_out <= "11010001"; -- 0xd1
                when "0001110010" => data_out <= "11010010"; -- 0xd2
                when "0001110011" => data_out <= "11010011"; -- 0xd3
                when "0001110100" => data_out <= "11010011"; -- 0xd3
                when "0001110101" => data_out <= "11010100"; -- 0xd4
                when "0001110110" => data_out <= "11010100"; -- 0xd4
                when "0001110111" => data_out <= "11010101"; -- 0xd5
                when "0001111000" => data_out <= "11010110"; -- 0xd6
                when "0001111001" => data_out <= "11010110"; -- 0xd6
                when "0001111010" => data_out <= "11010111"; -- 0xd7
                when "0001111011" => data_out <= "11010111"; -- 0xd7
                when "0001111100" => data_out <= "11011000"; -- 0xd8
                when "0001111101" => data_out <= "11011000"; -- 0xd8
                when "0001111110" => data_out <= "11011001"; -- 0xd9
                when "0001111111" => data_out <= "11011010"; -- 0xda
                when "0010000000" => data_out <= "11011010"; -- 0xda
                when "0010000001" => data_out <= "11011011"; -- 0xdb
                when "0010000010" => data_out <= "11011011"; -- 0xdb
                when "0010000011" => data_out <= "11011100"; -- 0xdc
                when "0010000100" => data_out <= "11011100"; -- 0xdc
                when "0010000101" => data_out <= "11011101"; -- 0xdd
                when "0010000110" => data_out <= "11011101"; -- 0xdd
                when "0010000111" => data_out <= "11011110"; -- 0xde
                when "0010001000" => data_out <= "11011110"; -- 0xde
                when "0010001001" => data_out <= "11011111"; -- 0xdf
                when "0010001010" => data_out <= "11011111"; -- 0xdf
                when "0010001011" => data_out <= "11100000"; -- 0xe0
                when "0010001100" => data_out <= "11100000"; -- 0xe0
                when "0010001101" => data_out <= "11100001"; -- 0xe1
                when "0010001110" => data_out <= "11100010"; -- 0xe2
                when "0010001111" => data_out <= "11100010"; -- 0xe2
                when "0010010000" => data_out <= "11100011"; -- 0xe3
                when "0010010001" => data_out <= "11100011"; -- 0xe3
                when "0010010010" => data_out <= "11100100"; -- 0xe4
                when "0010010011" => data_out <= "11100100"; -- 0xe4
                when "0010010100" => data_out <= "11100100"; -- 0xe4
                when "0010010101" => data_out <= "11100101"; -- 0xe5
                when "0010010110" => data_out <= "11100101"; -- 0xe5
                when "0010010111" => data_out <= "11100110"; -- 0xe6
                when "0010011000" => data_out <= "11100110"; -- 0xe6
                when "0010011001" => data_out <= "11100111"; -- 0xe7
                when "0010011010" => data_out <= "11100111"; -- 0xe7
                when "0010011011" => data_out <= "11101000"; -- 0xe8
                when "0010011100" => data_out <= "11101000"; -- 0xe8
                when "0010011101" => data_out <= "11101001"; -- 0xe9
                when "0010011110" => data_out <= "11101001"; -- 0xe9
                when "0010011111" => data_out <= "11101010"; -- 0xea
                when "0010100000" => data_out <= "11101010"; -- 0xea
                when "0010100001" => data_out <= "11101010"; -- 0xea
                when "0010100010" => data_out <= "11101011"; -- 0xeb
                when "0010100011" => data_out <= "11101011"; -- 0xeb
                when "0010100100" => data_out <= "11101100"; -- 0xec
                when "0010100101" => data_out <= "11101100"; -- 0xec
                when "0010100110" => data_out <= "11101101"; -- 0xed
                when "0010100111" => data_out <= "11101101"; -- 0xed
                when "0010101000" => data_out <= "11101101"; -- 0xed
                when "0010101001" => data_out <= "11101110"; -- 0xee
                when "0010101010" => data_out <= "11101110"; -- 0xee
                when "0010101011" => data_out <= "11101111"; -- 0xef
                when "0010101100" => data_out <= "11101111"; -- 0xef
                when "0010101101" => data_out <= "11101111"; -- 0xef
                when "0010101110" => data_out <= "11110000"; -- 0xf0
                when "0010101111" => data_out <= "11110000"; -- 0xf0
                when "0010110000" => data_out <= "11110000"; -- 0xf0
                when "0010110001" => data_out <= "11110001"; -- 0xf1
                when "0010110010" => data_out <= "11110001"; -- 0xf1
                when "0010110011" => data_out <= "11110010"; -- 0xf2
                when "0010110100" => data_out <= "11110010"; -- 0xf2
                when "0010110101" => data_out <= "11110010"; -- 0xf2
                when "0010110110" => data_out <= "11110011"; -- 0xf3
                when "0010110111" => data_out <= "11110011"; -- 0xf3
                when "0010111000" => data_out <= "11110011"; -- 0xf3
                when "0010111001" => data_out <= "11110100"; -- 0xf4
                when "0010111010" => data_out <= "11110100"; -- 0xf4
                when "0010111011" => data_out <= "11110100"; -- 0xf4
                when "0010111100" => data_out <= "11110101"; -- 0xf5
                when "0010111101" => data_out <= "11110101"; -- 0xf5
                when "0010111110" => data_out <= "11110101"; -- 0xf5
                when "0010111111" => data_out <= "11110110"; -- 0xf6
                when "0011000000" => data_out <= "11110110"; -- 0xf6
                when "0011000001" => data_out <= "11110110"; -- 0xf6
                when "0011000010" => data_out <= "11110110"; -- 0xf6
                when "0011000011" => data_out <= "11110111"; -- 0xf7
                when "0011000100" => data_out <= "11110111"; -- 0xf7
                when "0011000101" => data_out <= "11110111"; -- 0xf7
                when "0011000110" => data_out <= "11111000"; -- 0xf8
                when "0011000111" => data_out <= "11111000"; -- 0xf8
                when "0011001000" => data_out <= "11111000"; -- 0xf8
                when "0011001001" => data_out <= "11111000"; -- 0xf8
                when "0011001010" => data_out <= "11111001"; -- 0xf9
                when "0011001011" => data_out <= "11111001"; -- 0xf9
                when "0011001100" => data_out <= "11111001"; -- 0xf9
                when "0011001101" => data_out <= "11111001"; -- 0xf9
                when "0011001110" => data_out <= "11111010"; -- 0xfa
                when "0011001111" => data_out <= "11111010"; -- 0xfa
                when "0011010000" => data_out <= "11111010"; -- 0xfa
                when "0011010001" => data_out <= "11111010"; -- 0xfa
                when "0011010010" => data_out <= "11111010"; -- 0xfa
                when "0011010011" => data_out <= "11111011"; -- 0xfb
                when "0011010100" => data_out <= "11111011"; -- 0xfb
                when "0011010101" => data_out <= "11111011"; -- 0xfb
                when "0011010110" => data_out <= "11111011"; -- 0xfb
                when "0011010111" => data_out <= "11111100"; -- 0xfc
                when "0011011000" => data_out <= "11111100"; -- 0xfc
                when "0011011001" => data_out <= "11111100"; -- 0xfc
                when "0011011010" => data_out <= "11111100"; -- 0xfc
                when "0011011011" => data_out <= "11111100"; -- 0xfc
                when "0011011100" => data_out <= "11111100"; -- 0xfc
                when "0011011101" => data_out <= "11111101"; -- 0xfd
                when "0011011110" => data_out <= "11111101"; -- 0xfd
                when "0011011111" => data_out <= "11111101"; -- 0xfd
                when "0011100000" => data_out <= "11111101"; -- 0xfd
                when "0011100001" => data_out <= "11111101"; -- 0xfd
                when "0011100010" => data_out <= "11111101"; -- 0xfd
                when "0011100011" => data_out <= "11111110"; -- 0xfe
                when "0011100100" => data_out <= "11111110"; -- 0xfe
                when "0011100101" => data_out <= "11111110"; -- 0xfe
                when "0011100110" => data_out <= "11111110"; -- 0xfe
                when "0011100111" => data_out <= "11111110"; -- 0xfe
                when "0011101000" => data_out <= "11111110"; -- 0xfe
                when "0011101001" => data_out <= "11111110"; -- 0xfe
                when "0011101010" => data_out <= "11111110"; -- 0xfe
                when "0011101011" => data_out <= "11111110"; -- 0xfe
                when "0011101100" => data_out <= "11111111"; -- 0xff
                when "0011101101" => data_out <= "11111111"; -- 0xff
                when "0011101110" => data_out <= "11111111"; -- 0xff
                when "0011101111" => data_out <= "11111111"; -- 0xff
                when "0011110000" => data_out <= "11111111"; -- 0xff
                when "0011110001" => data_out <= "11111111"; -- 0xff
                when "0011110010" => data_out <= "11111111"; -- 0xff
                when "0011110011" => data_out <= "11111111"; -- 0xff
                when "0011110100" => data_out <= "11111111"; -- 0xff
                when "0011110101" => data_out <= "11111111"; -- 0xff
                when "0011110110" => data_out <= "11111111"; -- 0xff
                when "0011110111" => data_out <= "11111111"; -- 0xff
                when "0011111000" => data_out <= "11111111"; -- 0xff
                when "0011111001" => data_out <= "11111111"; -- 0xff
                when "0011111010" => data_out <= "11111111"; -- 0xff
                when "0011111011" => data_out <= "11111111"; -- 0xff
                when "0011111100" => data_out <= "11111111"; -- 0xff
                when "0011111101" => data_out <= "11111111"; -- 0xff
                when "0011111110" => data_out <= "11111111"; -- 0xff
                when "0011111111" => data_out <= "11111111"; -- 0xff
                when "0100000000" => data_out <= "11111111"; -- 0xff
                when "0100000001" => data_out <= "11111111"; -- 0xff
                when "0100000010" => data_out <= "11111111"; -- 0xff
                when "0100000011" => data_out <= "11111111"; -- 0xff
                when "0100000100" => data_out <= "11111111"; -- 0xff
                when "0100000101" => data_out <= "11111111"; -- 0xff
                when "0100000110" => data_out <= "11111111"; -- 0xff
                when "0100000111" => data_out <= "11111111"; -- 0xff
                when "0100001000" => data_out <= "11111111"; -- 0xff
                when "0100001001" => data_out <= "11111111"; -- 0xff
                when "0100001010" => data_out <= "11111111"; -- 0xff
                when "0100001011" => data_out <= "11111111"; -- 0xff
                when "0100001100" => data_out <= "11111111"; -- 0xff
                when "0100001101" => data_out <= "11111111"; -- 0xff
                when "0100001110" => data_out <= "11111111"; -- 0xff
                when "0100001111" => data_out <= "11111111"; -- 0xff
                when "0100010000" => data_out <= "11111111"; -- 0xff
                when "0100010001" => data_out <= "11111111"; -- 0xff
                when "0100010010" => data_out <= "11111111"; -- 0xff
                when "0100010011" => data_out <= "11111111"; -- 0xff
                when "0100010100" => data_out <= "11111111"; -- 0xff
                when "0100010101" => data_out <= "11111110"; -- 0xfe
                when "0100010110" => data_out <= "11111110"; -- 0xfe
                when "0100010111" => data_out <= "11111110"; -- 0xfe
                when "0100011000" => data_out <= "11111110"; -- 0xfe
                when "0100011001" => data_out <= "11111110"; -- 0xfe
                when "0100011010" => data_out <= "11111110"; -- 0xfe
                when "0100011011" => data_out <= "11111110"; -- 0xfe
                when "0100011100" => data_out <= "11111110"; -- 0xfe
                when "0100011101" => data_out <= "11111101"; -- 0xfd
                when "0100011110" => data_out <= "11111101"; -- 0xfd
                when "0100011111" => data_out <= "11111101"; -- 0xfd
                when "0100100000" => data_out <= "11111101"; -- 0xfd
                when "0100100001" => data_out <= "11111101"; -- 0xfd
                when "0100100010" => data_out <= "11111101"; -- 0xfd
                when "0100100011" => data_out <= "11111101"; -- 0xfd
                when "0100100100" => data_out <= "11111100"; -- 0xfc
                when "0100100101" => data_out <= "11111100"; -- 0xfc
                when "0100100110" => data_out <= "11111100"; -- 0xfc
                when "0100100111" => data_out <= "11111100"; -- 0xfc
                when "0100101000" => data_out <= "11111100"; -- 0xfc
                when "0100101001" => data_out <= "11111011"; -- 0xfb
                when "0100101010" => data_out <= "11111011"; -- 0xfb
                when "0100101011" => data_out <= "11111011"; -- 0xfb
                when "0100101100" => data_out <= "11111011"; -- 0xfb
                when "0100101101" => data_out <= "11111011"; -- 0xfb
                when "0100101110" => data_out <= "11111010"; -- 0xfa
                when "0100101111" => data_out <= "11111010"; -- 0xfa
                when "0100110000" => data_out <= "11111010"; -- 0xfa
                when "0100110001" => data_out <= "11111010"; -- 0xfa
                when "0100110010" => data_out <= "11111001"; -- 0xf9
                when "0100110011" => data_out <= "11111001"; -- 0xf9
                when "0100110100" => data_out <= "11111001"; -- 0xf9
                when "0100110101" => data_out <= "11111001"; -- 0xf9
                when "0100110110" => data_out <= "11111000"; -- 0xf8
                when "0100110111" => data_out <= "11111000"; -- 0xf8
                when "0100111000" => data_out <= "11111000"; -- 0xf8
                when "0100111001" => data_out <= "11111000"; -- 0xf8
                when "0100111010" => data_out <= "11110111"; -- 0xf7
                when "0100111011" => data_out <= "11110111"; -- 0xf7
                when "0100111100" => data_out <= "11110111"; -- 0xf7
                when "0100111101" => data_out <= "11110111"; -- 0xf7
                when "0100111110" => data_out <= "11110110"; -- 0xf6
                when "0100111111" => data_out <= "11110110"; -- 0xf6
                when "0101000000" => data_out <= "11110110"; -- 0xf6
                when "0101000001" => data_out <= "11110101"; -- 0xf5
                when "0101000010" => data_out <= "11110101"; -- 0xf5
                when "0101000011" => data_out <= "11110101"; -- 0xf5
                when "0101000100" => data_out <= "11110100"; -- 0xf4
                when "0101000101" => data_out <= "11110100"; -- 0xf4
                when "0101000110" => data_out <= "11110100"; -- 0xf4
                when "0101000111" => data_out <= "11110011"; -- 0xf3
                when "0101001000" => data_out <= "11110011"; -- 0xf3
                when "0101001001" => data_out <= "11110011"; -- 0xf3
                when "0101001010" => data_out <= "11110010"; -- 0xf2
                when "0101001011" => data_out <= "11110010"; -- 0xf2
                when "0101001100" => data_out <= "11110010"; -- 0xf2
                when "0101001101" => data_out <= "11110001"; -- 0xf1
                when "0101001110" => data_out <= "11110001"; -- 0xf1
                when "0101001111" => data_out <= "11110001"; -- 0xf1
                when "0101010000" => data_out <= "11110000"; -- 0xf0
                when "0101010001" => data_out <= "11110000"; -- 0xf0
                when "0101010010" => data_out <= "11110000"; -- 0xf0
                when "0101010011" => data_out <= "11101111"; -- 0xef
                when "0101010100" => data_out <= "11101111"; -- 0xef
                when "0101010101" => data_out <= "11101110"; -- 0xee
                when "0101010110" => data_out <= "11101110"; -- 0xee
                when "0101010111" => data_out <= "11101110"; -- 0xee
                when "0101011000" => data_out <= "11101101"; -- 0xed
                when "0101011001" => data_out <= "11101101"; -- 0xed
                when "0101011010" => data_out <= "11101100"; -- 0xec
                when "0101011011" => data_out <= "11101100"; -- 0xec
                when "0101011100" => data_out <= "11101011"; -- 0xeb
                when "0101011101" => data_out <= "11101011"; -- 0xeb
                when "0101011110" => data_out <= "11101011"; -- 0xeb
                when "0101011111" => data_out <= "11101010"; -- 0xea
                when "0101100000" => data_out <= "11101010"; -- 0xea
                when "0101100001" => data_out <= "11101001"; -- 0xe9
                when "0101100010" => data_out <= "11101001"; -- 0xe9
                when "0101100011" => data_out <= "11101000"; -- 0xe8
                when "0101100100" => data_out <= "11101000"; -- 0xe8
                when "0101100101" => data_out <= "11101000"; -- 0xe8
                when "0101100110" => data_out <= "11100111"; -- 0xe7
                when "0101100111" => data_out <= "11100111"; -- 0xe7
                when "0101101000" => data_out <= "11100110"; -- 0xe6
                when "0101101001" => data_out <= "11100110"; -- 0xe6
                when "0101101010" => data_out <= "11100101"; -- 0xe5
                when "0101101011" => data_out <= "11100101"; -- 0xe5
                when "0101101100" => data_out <= "11100100"; -- 0xe4
                when "0101101101" => data_out <= "11100100"; -- 0xe4
                when "0101101110" => data_out <= "11100011"; -- 0xe3
                when "0101101111" => data_out <= "11100011"; -- 0xe3
                when "0101110000" => data_out <= "11100010"; -- 0xe2
                when "0101110001" => data_out <= "11100010"; -- 0xe2
                when "0101110010" => data_out <= "11100001"; -- 0xe1
                when "0101110011" => data_out <= "11100001"; -- 0xe1
                when "0101110100" => data_out <= "11100000"; -- 0xe0
                when "0101110101" => data_out <= "11100000"; -- 0xe0
                when "0101110110" => data_out <= "11011111"; -- 0xdf
                when "0101110111" => data_out <= "11011111"; -- 0xdf
                when "0101111000" => data_out <= "11011110"; -- 0xde
                when "0101111001" => data_out <= "11011110"; -- 0xde
                when "0101111010" => data_out <= "11011101"; -- 0xdd
                when "0101111011" => data_out <= "11011101"; -- 0xdd
                when "0101111100" => data_out <= "11011100"; -- 0xdc
                when "0101111101" => data_out <= "11011011"; -- 0xdb
                when "0101111110" => data_out <= "11011011"; -- 0xdb
                when "0101111111" => data_out <= "11011010"; -- 0xda
                when "0110000000" => data_out <= "11011010"; -- 0xda
                when "0110000001" => data_out <= "11011001"; -- 0xd9
                when "0110000010" => data_out <= "11011001"; -- 0xd9
                when "0110000011" => data_out <= "11011000"; -- 0xd8
                when "0110000100" => data_out <= "11011000"; -- 0xd8
                when "0110000101" => data_out <= "11010111"; -- 0xd7
                when "0110000110" => data_out <= "11010110"; -- 0xd6
                when "0110000111" => data_out <= "11010110"; -- 0xd6
                when "0110001000" => data_out <= "11010101"; -- 0xd5
                when "0110001001" => data_out <= "11010101"; -- 0xd5
                when "0110001010" => data_out <= "11010100"; -- 0xd4
                when "0110001011" => data_out <= "11010011"; -- 0xd3
                when "0110001100" => data_out <= "11010011"; -- 0xd3
                when "0110001101" => data_out <= "11010010"; -- 0xd2
                when "0110001110" => data_out <= "11010010"; -- 0xd2
                when "0110001111" => data_out <= "11010001"; -- 0xd1
                when "0110010000" => data_out <= "11010000"; -- 0xd0
                when "0110010001" => data_out <= "11010000"; -- 0xd0
                when "0110010010" => data_out <= "11001111"; -- 0xcf
                when "0110010011" => data_out <= "11001111"; -- 0xcf
                when "0110010100" => data_out <= "11001110"; -- 0xce
                when "0110010101" => data_out <= "11001101"; -- 0xcd
                when "0110010110" => data_out <= "11001101"; -- 0xcd
                when "0110010111" => data_out <= "11001100"; -- 0xcc
                when "0110011000" => data_out <= "11001011"; -- 0xcb
                when "0110011001" => data_out <= "11001011"; -- 0xcb
                when "0110011010" => data_out <= "11001010"; -- 0xca
                when "0110011011" => data_out <= "11001010"; -- 0xca
                when "0110011100" => data_out <= "11001001"; -- 0xc9
                when "0110011101" => data_out <= "11001000"; -- 0xc8
                when "0110011110" => data_out <= "11001000"; -- 0xc8
                when "0110011111" => data_out <= "11000111"; -- 0xc7
                when "0110100000" => data_out <= "11000110"; -- 0xc6
                when "0110100001" => data_out <= "11000110"; -- 0xc6
                when "0110100010" => data_out <= "11000101"; -- 0xc5
                when "0110100011" => data_out <= "11000100"; -- 0xc4
                when "0110100100" => data_out <= "11000100"; -- 0xc4
                when "0110100101" => data_out <= "11000011"; -- 0xc3
                when "0110100110" => data_out <= "11000010"; -- 0xc2
                when "0110100111" => data_out <= "11000010"; -- 0xc2
                when "0110101000" => data_out <= "11000001"; -- 0xc1
                when "0110101001" => data_out <= "11000000"; -- 0xc0
                when "0110101010" => data_out <= "11000000"; -- 0xc0
                when "0110101011" => data_out <= "10111111"; -- 0xbf
                when "0110101100" => data_out <= "10111110"; -- 0xbe
                when "0110101101" => data_out <= "10111110"; -- 0xbe
                when "0110101110" => data_out <= "10111101"; -- 0xbd
                when "0110101111" => data_out <= "10111100"; -- 0xbc
                when "0110110000" => data_out <= "10111100"; -- 0xbc
                when "0110110001" => data_out <= "10111011"; -- 0xbb
                when "0110110010" => data_out <= "10111010"; -- 0xba
                when "0110110011" => data_out <= "10111001"; -- 0xb9
                when "0110110100" => data_out <= "10111001"; -- 0xb9
                when "0110110101" => data_out <= "10111000"; -- 0xb8
                when "0110110110" => data_out <= "10110111"; -- 0xb7
                when "0110110111" => data_out <= "10110111"; -- 0xb7
                when "0110111000" => data_out <= "10110110"; -- 0xb6
                when "0110111001" => data_out <= "10110101"; -- 0xb5
                when "0110111010" => data_out <= "10110100"; -- 0xb4
                when "0110111011" => data_out <= "10110100"; -- 0xb4
                when "0110111100" => data_out <= "10110011"; -- 0xb3
                when "0110111101" => data_out <= "10110010"; -- 0xb2
                when "0110111110" => data_out <= "10110010"; -- 0xb2
                when "0110111111" => data_out <= "10110001"; -- 0xb1
                when "0111000000" => data_out <= "10110000"; -- 0xb0
                when "0111000001" => data_out <= "10101111"; -- 0xaf
                when "0111000010" => data_out <= "10101111"; -- 0xaf
                when "0111000011" => data_out <= "10101110"; -- 0xae
                when "0111000100" => data_out <= "10101101"; -- 0xad
                when "0111000101" => data_out <= "10101101"; -- 0xad
                when "0111000110" => data_out <= "10101100"; -- 0xac
                when "0111000111" => data_out <= "10101011"; -- 0xab
                when "0111001000" => data_out <= "10101010"; -- 0xaa
                when "0111001001" => data_out <= "10101010"; -- 0xaa
                when "0111001010" => data_out <= "10101001"; -- 0xa9
                when "0111001011" => data_out <= "10101000"; -- 0xa8
                when "0111001100" => data_out <= "10100111"; -- 0xa7
                when "0111001101" => data_out <= "10100111"; -- 0xa7
                when "0111001110" => data_out <= "10100110"; -- 0xa6
                when "0111001111" => data_out <= "10100101"; -- 0xa5
                when "0111010000" => data_out <= "10100100"; -- 0xa4
                when "0111010001" => data_out <= "10100100"; -- 0xa4
                when "0111010010" => data_out <= "10100011"; -- 0xa3
                when "0111010011" => data_out <= "10100010"; -- 0xa2
                when "0111010100" => data_out <= "10100001"; -- 0xa1
                when "0111010101" => data_out <= "10100001"; -- 0xa1
                when "0111010110" => data_out <= "10100000"; -- 0xa0
                when "0111010111" => data_out <= "10011111"; -- 0x9f
                when "0111011000" => data_out <= "10011110"; -- 0x9e
                when "0111011001" => data_out <= "10011101"; -- 0x9d
                when "0111011010" => data_out <= "10011101"; -- 0x9d
                when "0111011011" => data_out <= "10011100"; -- 0x9c
                when "0111011100" => data_out <= "10011011"; -- 0x9b
                when "0111011101" => data_out <= "10011010"; -- 0x9a
                when "0111011110" => data_out <= "10011010"; -- 0x9a
                when "0111011111" => data_out <= "10011001"; -- 0x99
                when "0111100000" => data_out <= "10011000"; -- 0x98
                when "0111100001" => data_out <= "10010111"; -- 0x97
                when "0111100010" => data_out <= "10010111"; -- 0x97
                when "0111100011" => data_out <= "10010110"; -- 0x96
                when "0111100100" => data_out <= "10010101"; -- 0x95
                when "0111100101" => data_out <= "10010100"; -- 0x94
                when "0111100110" => data_out <= "10010011"; -- 0x93
                when "0111100111" => data_out <= "10010011"; -- 0x93
                when "0111101000" => data_out <= "10010010"; -- 0x92
                when "0111101001" => data_out <= "10010001"; -- 0x91
                when "0111101010" => data_out <= "10010000"; -- 0x90
                when "0111101011" => data_out <= "10010000"; -- 0x90
                when "0111101100" => data_out <= "10001111"; -- 0x8f
                when "0111101101" => data_out <= "10001110"; -- 0x8e
                when "0111101110" => data_out <= "10001101"; -- 0x8d
                when "0111101111" => data_out <= "10001100"; -- 0x8c
                when "0111110000" => data_out <= "10001100"; -- 0x8c
                when "0111110001" => data_out <= "10001011"; -- 0x8b
                when "0111110010" => data_out <= "10001010"; -- 0x8a
                when "0111110011" => data_out <= "10001001"; -- 0x89
                when "0111110100" => data_out <= "10001001"; -- 0x89
                when "0111110101" => data_out <= "10001000"; -- 0x88
                when "0111110110" => data_out <= "10000111"; -- 0x87
                when "0111110111" => data_out <= "10000110"; -- 0x86
                when "0111111000" => data_out <= "10000101"; -- 0x85
                when "0111111001" => data_out <= "10000101"; -- 0x85
                when "0111111010" => data_out <= "10000100"; -- 0x84
                when "0111111011" => data_out <= "10000011"; -- 0x83
                when "0111111100" => data_out <= "10000010"; -- 0x82
                when "0111111101" => data_out <= "10000001"; -- 0x81
                when "0111111110" => data_out <= "10000001"; -- 0x81
                when "0111111111" => data_out <= "10000000"; -- 0x80
                when "1000000000" => data_out <= "01111111"; -- 0x7f
                when "1000000001" => data_out <= "01111110"; -- 0x7e
                when "1000000010" => data_out <= "01111110"; -- 0x7e
                when "1000000011" => data_out <= "01111101"; -- 0x7d
                when "1000000100" => data_out <= "01111100"; -- 0x7c
                when "1000000101" => data_out <= "01111011"; -- 0x7b
                when "1000000110" => data_out <= "01111010"; -- 0x7a
                when "1000000111" => data_out <= "01111010"; -- 0x7a
                when "1000001000" => data_out <= "01111001"; -- 0x79
                when "1000001001" => data_out <= "01111000"; -- 0x78
                when "1000001010" => data_out <= "01110111"; -- 0x77
                when "1000001011" => data_out <= "01110110"; -- 0x76
                when "1000001100" => data_out <= "01110110"; -- 0x76
                when "1000001101" => data_out <= "01110101"; -- 0x75
                when "1000001110" => data_out <= "01110100"; -- 0x74
                when "1000001111" => data_out <= "01110011"; -- 0x73
                when "1000010000" => data_out <= "01110011"; -- 0x73
                when "1000010001" => data_out <= "01110010"; -- 0x72
                when "1000010010" => data_out <= "01110001"; -- 0x71
                when "1000010011" => data_out <= "01110000"; -- 0x70
                when "1000010100" => data_out <= "01101111"; -- 0x6f
                when "1000010101" => data_out <= "01101111"; -- 0x6f
                when "1000010110" => data_out <= "01101110"; -- 0x6e
                when "1000010111" => data_out <= "01101101"; -- 0x6d
                when "1000011000" => data_out <= "01101100"; -- 0x6c
                when "1000011001" => data_out <= "01101100"; -- 0x6c
                when "1000011010" => data_out <= "01101011"; -- 0x6b
                when "1000011011" => data_out <= "01101010"; -- 0x6a
                when "1000011100" => data_out <= "01101001"; -- 0x69
                when "1000011101" => data_out <= "01101000"; -- 0x68
                when "1000011110" => data_out <= "01101000"; -- 0x68
                when "1000011111" => data_out <= "01100111"; -- 0x67
                when "1000100000" => data_out <= "01100110"; -- 0x66
                when "1000100001" => data_out <= "01100101"; -- 0x65
                when "1000100010" => data_out <= "01100101"; -- 0x65
                when "1000100011" => data_out <= "01100100"; -- 0x64
                when "1000100100" => data_out <= "01100011"; -- 0x63
                when "1000100101" => data_out <= "01100010"; -- 0x62
                when "1000100110" => data_out <= "01100010"; -- 0x62
                when "1000100111" => data_out <= "01100001"; -- 0x61
                when "1000101000" => data_out <= "01100000"; -- 0x60
                when "1000101001" => data_out <= "01011111"; -- 0x5f
                when "1000101010" => data_out <= "01011110"; -- 0x5e
                when "1000101011" => data_out <= "01011110"; -- 0x5e
                when "1000101100" => data_out <= "01011101"; -- 0x5d
                when "1000101101" => data_out <= "01011100"; -- 0x5c
                when "1000101110" => data_out <= "01011011"; -- 0x5b
                when "1000101111" => data_out <= "01011011"; -- 0x5b
                when "1000110000" => data_out <= "01011010"; -- 0x5a
                when "1000110001" => data_out <= "01011001"; -- 0x59
                when "1000110010" => data_out <= "01011000"; -- 0x58
                when "1000110011" => data_out <= "01011000"; -- 0x58
                when "1000110100" => data_out <= "01010111"; -- 0x57
                when "1000110101" => data_out <= "01010110"; -- 0x56
                when "1000110110" => data_out <= "01010101"; -- 0x55
                when "1000110111" => data_out <= "01010101"; -- 0x55
                when "1000111000" => data_out <= "01010100"; -- 0x54
                when "1000111001" => data_out <= "01010011"; -- 0x53
                when "1000111010" => data_out <= "01010010"; -- 0x52
                when "1000111011" => data_out <= "01010010"; -- 0x52
                when "1000111100" => data_out <= "01010001"; -- 0x51
                when "1000111101" => data_out <= "01010000"; -- 0x50
                when "1000111110" => data_out <= "01010000"; -- 0x50
                when "1000111111" => data_out <= "01001111"; -- 0x4f
                when "1001000000" => data_out <= "01001110"; -- 0x4e
                when "1001000001" => data_out <= "01001101"; -- 0x4d
                when "1001000010" => data_out <= "01001101"; -- 0x4d
                when "1001000011" => data_out <= "01001100"; -- 0x4c
                when "1001000100" => data_out <= "01001011"; -- 0x4b
                when "1001000101" => data_out <= "01001011"; -- 0x4b
                when "1001000110" => data_out <= "01001010"; -- 0x4a
                when "1001000111" => data_out <= "01001001"; -- 0x49
                when "1001001000" => data_out <= "01001000"; -- 0x48
                when "1001001001" => data_out <= "01001000"; -- 0x48
                when "1001001010" => data_out <= "01000111"; -- 0x47
                when "1001001011" => data_out <= "01000110"; -- 0x46
                when "1001001100" => data_out <= "01000110"; -- 0x46
                when "1001001101" => data_out <= "01000101"; -- 0x45
                when "1001001110" => data_out <= "01000100"; -- 0x44
                when "1001001111" => data_out <= "01000011"; -- 0x43
                when "1001010000" => data_out <= "01000011"; -- 0x43
                when "1001010001" => data_out <= "01000010"; -- 0x42
                when "1001010010" => data_out <= "01000001"; -- 0x41
                when "1001010011" => data_out <= "01000001"; -- 0x41
                when "1001010100" => data_out <= "01000000"; -- 0x40
                when "1001010101" => data_out <= "00111111"; -- 0x3f
                when "1001010110" => data_out <= "00111111"; -- 0x3f
                when "1001010111" => data_out <= "00111110"; -- 0x3e
                when "1001011000" => data_out <= "00111101"; -- 0x3d
                when "1001011001" => data_out <= "00111101"; -- 0x3d
                when "1001011010" => data_out <= "00111100"; -- 0x3c
                when "1001011011" => data_out <= "00111011"; -- 0x3b
                when "1001011100" => data_out <= "00111011"; -- 0x3b
                when "1001011101" => data_out <= "00111010"; -- 0x3a
                when "1001011110" => data_out <= "00111001"; -- 0x39
                when "1001011111" => data_out <= "00111001"; -- 0x39
                when "1001100000" => data_out <= "00111000"; -- 0x38
                when "1001100001" => data_out <= "00110111"; -- 0x37
                when "1001100010" => data_out <= "00110111"; -- 0x37
                when "1001100011" => data_out <= "00110110"; -- 0x36
                when "1001100100" => data_out <= "00110101"; -- 0x35
                when "1001100101" => data_out <= "00110101"; -- 0x35
                when "1001100110" => data_out <= "00110100"; -- 0x34
                when "1001100111" => data_out <= "00110100"; -- 0x34
                when "1001101000" => data_out <= "00110011"; -- 0x33
                when "1001101001" => data_out <= "00110010"; -- 0x32
                when "1001101010" => data_out <= "00110010"; -- 0x32
                when "1001101011" => data_out <= "00110001"; -- 0x31
                when "1001101100" => data_out <= "00110000"; -- 0x30
                when "1001101101" => data_out <= "00110000"; -- 0x30
                when "1001101110" => data_out <= "00101111"; -- 0x2f
                when "1001101111" => data_out <= "00101111"; -- 0x2f
                when "1001110000" => data_out <= "00101110"; -- 0x2e
                when "1001110001" => data_out <= "00101101"; -- 0x2d
                when "1001110010" => data_out <= "00101101"; -- 0x2d
                when "1001110011" => data_out <= "00101100"; -- 0x2c
                when "1001110100" => data_out <= "00101100"; -- 0x2c
                when "1001110101" => data_out <= "00101011"; -- 0x2b
                when "1001110110" => data_out <= "00101010"; -- 0x2a
                when "1001110111" => data_out <= "00101010"; -- 0x2a
                when "1001111000" => data_out <= "00101001"; -- 0x29
                when "1001111001" => data_out <= "00101001"; -- 0x29
                when "1001111010" => data_out <= "00101000"; -- 0x28
                when "1001111011" => data_out <= "00100111"; -- 0x27
                when "1001111100" => data_out <= "00100111"; -- 0x27
                when "1001111101" => data_out <= "00100110"; -- 0x26
                when "1001111110" => data_out <= "00100110"; -- 0x26
                when "1001111111" => data_out <= "00100101"; -- 0x25
                when "1010000000" => data_out <= "00100101"; -- 0x25
                when "1010000001" => data_out <= "00100100"; -- 0x24
                when "1010000010" => data_out <= "00100100"; -- 0x24
                when "1010000011" => data_out <= "00100011"; -- 0x23
                when "1010000100" => data_out <= "00100010"; -- 0x22
                when "1010000101" => data_out <= "00100010"; -- 0x22
                when "1010000110" => data_out <= "00100001"; -- 0x21
                when "1010000111" => data_out <= "00100001"; -- 0x21
                when "1010001000" => data_out <= "00100000"; -- 0x20
                when "1010001001" => data_out <= "00100000"; -- 0x20
                when "1010001010" => data_out <= "00011111"; -- 0x1f
                when "1010001011" => data_out <= "00011111"; -- 0x1f
                when "1010001100" => data_out <= "00011110"; -- 0x1e
                when "1010001101" => data_out <= "00011110"; -- 0x1e
                when "1010001110" => data_out <= "00011101"; -- 0x1d
                when "1010001111" => data_out <= "00011101"; -- 0x1d
                when "1010010000" => data_out <= "00011100"; -- 0x1c
                when "1010010001" => data_out <= "00011100"; -- 0x1c
                when "1010010010" => data_out <= "00011011"; -- 0x1b
                when "1010010011" => data_out <= "00011011"; -- 0x1b
                when "1010010100" => data_out <= "00011010"; -- 0x1a
                when "1010010101" => data_out <= "00011010"; -- 0x1a
                when "1010010110" => data_out <= "00011001"; -- 0x19
                when "1010010111" => data_out <= "00011001"; -- 0x19
                when "1010011000" => data_out <= "00011000"; -- 0x18
                when "1010011001" => data_out <= "00011000"; -- 0x18
                when "1010011010" => data_out <= "00010111"; -- 0x17
                when "1010011011" => data_out <= "00010111"; -- 0x17
                when "1010011100" => data_out <= "00010111"; -- 0x17
                when "1010011101" => data_out <= "00010110"; -- 0x16
                when "1010011110" => data_out <= "00010110"; -- 0x16
                when "1010011111" => data_out <= "00010101"; -- 0x15
                when "1010100000" => data_out <= "00010101"; -- 0x15
                when "1010100001" => data_out <= "00010100"; -- 0x14
                when "1010100010" => data_out <= "00010100"; -- 0x14
                when "1010100011" => data_out <= "00010100"; -- 0x14
                when "1010100100" => data_out <= "00010011"; -- 0x13
                when "1010100101" => data_out <= "00010011"; -- 0x13
                when "1010100110" => data_out <= "00010010"; -- 0x12
                when "1010100111" => data_out <= "00010010"; -- 0x12
                when "1010101000" => data_out <= "00010001"; -- 0x11
                when "1010101001" => data_out <= "00010001"; -- 0x11
                when "1010101010" => data_out <= "00010001"; -- 0x11
                when "1010101011" => data_out <= "00010000"; -- 0x10
                when "1010101100" => data_out <= "00010000"; -- 0x10
                when "1010101101" => data_out <= "00001111"; -- 0xf
                when "1010101110" => data_out <= "00001111"; -- 0xf
                when "1010101111" => data_out <= "00001111"; -- 0xf
                when "1010110000" => data_out <= "00001110"; -- 0xe
                when "1010110001" => data_out <= "00001110"; -- 0xe
                when "1010110010" => data_out <= "00001110"; -- 0xe
                when "1010110011" => data_out <= "00001101"; -- 0xd
                when "1010110100" => data_out <= "00001101"; -- 0xd
                when "1010110101" => data_out <= "00001101"; -- 0xd
                when "1010110110" => data_out <= "00001100"; -- 0xc
                when "1010110111" => data_out <= "00001100"; -- 0xc
                when "1010111000" => data_out <= "00001100"; -- 0xc
                when "1010111001" => data_out <= "00001011"; -- 0xb
                when "1010111010" => data_out <= "00001011"; -- 0xb
                when "1010111011" => data_out <= "00001011"; -- 0xb
                when "1010111100" => data_out <= "00001010"; -- 0xa
                when "1010111101" => data_out <= "00001010"; -- 0xa
                when "1010111110" => data_out <= "00001010"; -- 0xa
                when "1010111111" => data_out <= "00001001"; -- 0x9
                when "1011000000" => data_out <= "00001001"; -- 0x9
                when "1011000001" => data_out <= "00001001"; -- 0x9
                when "1011000010" => data_out <= "00001000"; -- 0x8
                when "1011000011" => data_out <= "00001000"; -- 0x8
                when "1011000100" => data_out <= "00001000"; -- 0x8
                when "1011000101" => data_out <= "00001000"; -- 0x8
                when "1011000110" => data_out <= "00000111"; -- 0x7
                when "1011000111" => data_out <= "00000111"; -- 0x7
                when "1011001000" => data_out <= "00000111"; -- 0x7
                when "1011001001" => data_out <= "00000111"; -- 0x7
                when "1011001010" => data_out <= "00000110"; -- 0x6
                when "1011001011" => data_out <= "00000110"; -- 0x6
                when "1011001100" => data_out <= "00000110"; -- 0x6
                when "1011001101" => data_out <= "00000110"; -- 0x6
                when "1011001110" => data_out <= "00000101"; -- 0x5
                when "1011001111" => data_out <= "00000101"; -- 0x5
                when "1011010000" => data_out <= "00000101"; -- 0x5
                when "1011010001" => data_out <= "00000101"; -- 0x5
                when "1011010010" => data_out <= "00000100"; -- 0x4
                when "1011010011" => data_out <= "00000100"; -- 0x4
                when "1011010100" => data_out <= "00000100"; -- 0x4
                when "1011010101" => data_out <= "00000100"; -- 0x4
                when "1011010110" => data_out <= "00000100"; -- 0x4
                when "1011010111" => data_out <= "00000011"; -- 0x3
                when "1011011000" => data_out <= "00000011"; -- 0x3
                when "1011011001" => data_out <= "00000011"; -- 0x3
                when "1011011010" => data_out <= "00000011"; -- 0x3
                when "1011011011" => data_out <= "00000011"; -- 0x3
                when "1011011100" => data_out <= "00000010"; -- 0x2
                when "1011011101" => data_out <= "00000010"; -- 0x2
                when "1011011110" => data_out <= "00000010"; -- 0x2
                when "1011011111" => data_out <= "00000010"; -- 0x2
                when "1011100000" => data_out <= "00000010"; -- 0x2
                when "1011100001" => data_out <= "00000010"; -- 0x2
                when "1011100010" => data_out <= "00000010"; -- 0x2
                when "1011100011" => data_out <= "00000001"; -- 0x1
                when "1011100100" => data_out <= "00000001"; -- 0x1
                when "1011100101" => data_out <= "00000001"; -- 0x1
                when "1011100110" => data_out <= "00000001"; -- 0x1
                when "1011100111" => data_out <= "00000001"; -- 0x1
                when "1011101000" => data_out <= "00000001"; -- 0x1
                when "1011101001" => data_out <= "00000001"; -- 0x1
                when "1011101010" => data_out <= "00000001"; -- 0x1
                when "1011101011" => data_out <= "00000000"; -- 0x0
                when "1011101100" => data_out <= "00000000"; -- 0x0
                when "1011101101" => data_out <= "00000000"; -- 0x0
                when "1011101110" => data_out <= "00000000"; -- 0x0
                when "1011101111" => data_out <= "00000000"; -- 0x0
                when "1011110000" => data_out <= "00000000"; -- 0x0
                when "1011110001" => data_out <= "00000000"; -- 0x0
                when "1011110010" => data_out <= "00000000"; -- 0x0
                when "1011110011" => data_out <= "00000000"; -- 0x0
                when "1011110100" => data_out <= "00000000"; -- 0x0
                when "1011110101" => data_out <= "00000000"; -- 0x0
                when "1011110110" => data_out <= "00000000"; -- 0x0
                when "1011110111" => data_out <= "00000000"; -- 0x0
                when "1011111000" => data_out <= "00000000"; -- 0x0
                when "1011111001" => data_out <= "00000000"; -- 0x0
                when "1011111010" => data_out <= "00000000"; -- 0x0
                when "1011111011" => data_out <= "00000000"; -- 0x0
                when "1011111100" => data_out <= "00000000"; -- 0x0
                when "1011111101" => data_out <= "00000000"; -- 0x0
                when "1011111110" => data_out <= "00000000"; -- 0x0
                when "1011111111" => data_out <= "00000000"; -- 0x0
                when "1100000000" => data_out <= "00000000"; -- 0x0
                when "1100000001" => data_out <= "00000000"; -- 0x0
                when "1100000010" => data_out <= "00000000"; -- 0x0
                when "1100000011" => data_out <= "00000000"; -- 0x0
                when "1100000100" => data_out <= "00000000"; -- 0x0
                when "1100000101" => data_out <= "00000000"; -- 0x0
                when "1100000110" => data_out <= "00000000"; -- 0x0
                when "1100000111" => data_out <= "00000000"; -- 0x0
                when "1100001000" => data_out <= "00000000"; -- 0x0
                when "1100001001" => data_out <= "00000000"; -- 0x0
                when "1100001010" => data_out <= "00000000"; -- 0x0
                when "1100001011" => data_out <= "00000000"; -- 0x0
                when "1100001100" => data_out <= "00000000"; -- 0x0
                when "1100001101" => data_out <= "00000000"; -- 0x0
                when "1100001110" => data_out <= "00000000"; -- 0x0
                when "1100001111" => data_out <= "00000000"; -- 0x0
                when "1100010000" => data_out <= "00000000"; -- 0x0
                when "1100010001" => data_out <= "00000000"; -- 0x0
                when "1100010010" => data_out <= "00000000"; -- 0x0
                when "1100010011" => data_out <= "00000000"; -- 0x0
                when "1100010100" => data_out <= "00000001"; -- 0x1
                when "1100010101" => data_out <= "00000001"; -- 0x1
                when "1100010110" => data_out <= "00000001"; -- 0x1
                when "1100010111" => data_out <= "00000001"; -- 0x1
                when "1100011000" => data_out <= "00000001"; -- 0x1
                when "1100011001" => data_out <= "00000001"; -- 0x1
                when "1100011010" => data_out <= "00000001"; -- 0x1
                when "1100011011" => data_out <= "00000001"; -- 0x1
                when "1100011100" => data_out <= "00000001"; -- 0x1
                when "1100011101" => data_out <= "00000010"; -- 0x2
                when "1100011110" => data_out <= "00000010"; -- 0x2
                when "1100011111" => data_out <= "00000010"; -- 0x2
                when "1100100000" => data_out <= "00000010"; -- 0x2
                when "1100100001" => data_out <= "00000010"; -- 0x2
                when "1100100010" => data_out <= "00000010"; -- 0x2
                when "1100100011" => data_out <= "00000011"; -- 0x3
                when "1100100100" => data_out <= "00000011"; -- 0x3
                when "1100100101" => data_out <= "00000011"; -- 0x3
                when "1100100110" => data_out <= "00000011"; -- 0x3
                when "1100100111" => data_out <= "00000011"; -- 0x3
                when "1100101000" => data_out <= "00000011"; -- 0x3
                when "1100101001" => data_out <= "00000100"; -- 0x4
                when "1100101010" => data_out <= "00000100"; -- 0x4
                when "1100101011" => data_out <= "00000100"; -- 0x4
                when "1100101100" => data_out <= "00000100"; -- 0x4
                when "1100101101" => data_out <= "00000101"; -- 0x5
                when "1100101110" => data_out <= "00000101"; -- 0x5
                when "1100101111" => data_out <= "00000101"; -- 0x5
                when "1100110000" => data_out <= "00000101"; -- 0x5
                when "1100110001" => data_out <= "00000101"; -- 0x5
                when "1100110010" => data_out <= "00000110"; -- 0x6
                when "1100110011" => data_out <= "00000110"; -- 0x6
                when "1100110100" => data_out <= "00000110"; -- 0x6
                when "1100110101" => data_out <= "00000110"; -- 0x6
                when "1100110110" => data_out <= "00000111"; -- 0x7
                when "1100110111" => data_out <= "00000111"; -- 0x7
                when "1100111000" => data_out <= "00000111"; -- 0x7
                when "1100111001" => data_out <= "00000111"; -- 0x7
                when "1100111010" => data_out <= "00001000"; -- 0x8
                when "1100111011" => data_out <= "00001000"; -- 0x8
                when "1100111100" => data_out <= "00001000"; -- 0x8
                when "1100111101" => data_out <= "00001001"; -- 0x9
                when "1100111110" => data_out <= "00001001"; -- 0x9
                when "1100111111" => data_out <= "00001001"; -- 0x9
                when "1101000000" => data_out <= "00001001"; -- 0x9
                when "1101000001" => data_out <= "00001010"; -- 0xa
                when "1101000010" => data_out <= "00001010"; -- 0xa
                when "1101000011" => data_out <= "00001010"; -- 0xa
                when "1101000100" => data_out <= "00001011"; -- 0xb
                when "1101000101" => data_out <= "00001011"; -- 0xb
                when "1101000110" => data_out <= "00001011"; -- 0xb
                when "1101000111" => data_out <= "00001100"; -- 0xc
                when "1101001000" => data_out <= "00001100"; -- 0xc
                when "1101001001" => data_out <= "00001100"; -- 0xc
                when "1101001010" => data_out <= "00001101"; -- 0xd
                when "1101001011" => data_out <= "00001101"; -- 0xd
                when "1101001100" => data_out <= "00001101"; -- 0xd
                when "1101001101" => data_out <= "00001110"; -- 0xe
                when "1101001110" => data_out <= "00001110"; -- 0xe
                when "1101001111" => data_out <= "00001111"; -- 0xf
                when "1101010000" => data_out <= "00001111"; -- 0xf
                when "1101010001" => data_out <= "00001111"; -- 0xf
                when "1101010010" => data_out <= "00010000"; -- 0x10
                when "1101010011" => data_out <= "00010000"; -- 0x10
                when "1101010100" => data_out <= "00010000"; -- 0x10
                when "1101010101" => data_out <= "00010001"; -- 0x11
                when "1101010110" => data_out <= "00010001"; -- 0x11
                when "1101010111" => data_out <= "00010010"; -- 0x12
                when "1101011000" => data_out <= "00010010"; -- 0x12
                when "1101011001" => data_out <= "00010010"; -- 0x12
                when "1101011010" => data_out <= "00010011"; -- 0x13
                when "1101011011" => data_out <= "00010011"; -- 0x13
                when "1101011100" => data_out <= "00010100"; -- 0x14
                when "1101011101" => data_out <= "00010100"; -- 0x14
                when "1101011110" => data_out <= "00010101"; -- 0x15
                when "1101011111" => data_out <= "00010101"; -- 0x15
                when "1101100000" => data_out <= "00010101"; -- 0x15
                when "1101100001" => data_out <= "00010110"; -- 0x16
                when "1101100010" => data_out <= "00010110"; -- 0x16
                when "1101100011" => data_out <= "00010111"; -- 0x17
                when "1101100100" => data_out <= "00010111"; -- 0x17
                when "1101100101" => data_out <= "00011000"; -- 0x18
                when "1101100110" => data_out <= "00011000"; -- 0x18
                when "1101100111" => data_out <= "00011001"; -- 0x19
                when "1101101000" => data_out <= "00011001"; -- 0x19
                when "1101101001" => data_out <= "00011010"; -- 0x1a
                when "1101101010" => data_out <= "00011010"; -- 0x1a
                when "1101101011" => data_out <= "00011011"; -- 0x1b
                when "1101101100" => data_out <= "00011011"; -- 0x1b
                when "1101101101" => data_out <= "00011011"; -- 0x1b
                when "1101101110" => data_out <= "00011100"; -- 0x1c
                when "1101101111" => data_out <= "00011100"; -- 0x1c
                when "1101110000" => data_out <= "00011101"; -- 0x1d
                when "1101110001" => data_out <= "00011101"; -- 0x1d
                when "1101110010" => data_out <= "00011110"; -- 0x1e
                when "1101110011" => data_out <= "00011111"; -- 0x1f
                when "1101110100" => data_out <= "00011111"; -- 0x1f
                when "1101110101" => data_out <= "00100000"; -- 0x20
                when "1101110110" => data_out <= "00100000"; -- 0x20
                when "1101110111" => data_out <= "00100001"; -- 0x21
                when "1101111000" => data_out <= "00100001"; -- 0x21
                when "1101111001" => data_out <= "00100010"; -- 0x22
                when "1101111010" => data_out <= "00100010"; -- 0x22
                when "1101111011" => data_out <= "00100011"; -- 0x23
                when "1101111100" => data_out <= "00100011"; -- 0x23
                when "1101111101" => data_out <= "00100100"; -- 0x24
                when "1101111110" => data_out <= "00100100"; -- 0x24
                when "1101111111" => data_out <= "00100101"; -- 0x25
                when "1110000000" => data_out <= "00100101"; -- 0x25
                when "1110000001" => data_out <= "00100110"; -- 0x26
                when "1110000010" => data_out <= "00100111"; -- 0x27
                when "1110000011" => data_out <= "00100111"; -- 0x27
                when "1110000100" => data_out <= "00101000"; -- 0x28
                when "1110000101" => data_out <= "00101000"; -- 0x28
                when "1110000110" => data_out <= "00101001"; -- 0x29
                when "1110000111" => data_out <= "00101001"; -- 0x29
                when "1110001000" => data_out <= "00101010"; -- 0x2a
                when "1110001001" => data_out <= "00101011"; -- 0x2b
                when "1110001010" => data_out <= "00101011"; -- 0x2b
                when "1110001011" => data_out <= "00101100"; -- 0x2c
                when "1110001100" => data_out <= "00101100"; -- 0x2c
                when "1110001101" => data_out <= "00101101"; -- 0x2d
                when "1110001110" => data_out <= "00101110"; -- 0x2e
                when "1110001111" => data_out <= "00101110"; -- 0x2e
                when "1110010000" => data_out <= "00101111"; -- 0x2f
                when "1110010001" => data_out <= "00101111"; -- 0x2f
                when "1110010010" => data_out <= "00110000"; -- 0x30
                when "1110010011" => data_out <= "00110001"; -- 0x31
                when "1110010100" => data_out <= "00110001"; -- 0x31
                when "1110010101" => data_out <= "00110010"; -- 0x32
                when "1110010110" => data_out <= "00110011"; -- 0x33
                when "1110010111" => data_out <= "00110011"; -- 0x33
                when "1110011000" => data_out <= "00110100"; -- 0x34
                when "1110011001" => data_out <= "00110100"; -- 0x34
                when "1110011010" => data_out <= "00110101"; -- 0x35
                when "1110011011" => data_out <= "00110110"; -- 0x36
                when "1110011100" => data_out <= "00110110"; -- 0x36
                when "1110011101" => data_out <= "00110111"; -- 0x37
                when "1110011110" => data_out <= "00111000"; -- 0x38
                when "1110011111" => data_out <= "00111000"; -- 0x38
                when "1110100000" => data_out <= "00111001"; -- 0x39
                when "1110100001" => data_out <= "00111010"; -- 0x3a
                when "1110100010" => data_out <= "00111010"; -- 0x3a
                when "1110100011" => data_out <= "00111011"; -- 0x3b
                when "1110100100" => data_out <= "00111100"; -- 0x3c
                when "1110100101" => data_out <= "00111100"; -- 0x3c
                when "1110100110" => data_out <= "00111101"; -- 0x3d
                when "1110100111" => data_out <= "00111110"; -- 0x3e
                when "1110101000" => data_out <= "00111110"; -- 0x3e
                when "1110101001" => data_out <= "00111111"; -- 0x3f
                when "1110101010" => data_out <= "01000000"; -- 0x40
                when "1110101011" => data_out <= "01000000"; -- 0x40
                when "1110101100" => data_out <= "01000001"; -- 0x41
                when "1110101101" => data_out <= "01000010"; -- 0x42
                when "1110101110" => data_out <= "01000010"; -- 0x42
                when "1110101111" => data_out <= "01000011"; -- 0x43
                when "1110110000" => data_out <= "01000100"; -- 0x44
                when "1110110001" => data_out <= "01000100"; -- 0x44
                when "1110110010" => data_out <= "01000101"; -- 0x45
                when "1110110011" => data_out <= "01000110"; -- 0x46
                when "1110110100" => data_out <= "01000111"; -- 0x47
                when "1110110101" => data_out <= "01000111"; -- 0x47
                when "1110110110" => data_out <= "01001000"; -- 0x48
                when "1110110111" => data_out <= "01001001"; -- 0x49
                when "1110111000" => data_out <= "01001001"; -- 0x49
                when "1110111001" => data_out <= "01001010"; -- 0x4a
                when "1110111010" => data_out <= "01001011"; -- 0x4b
                when "1110111011" => data_out <= "01001100"; -- 0x4c
                when "1110111100" => data_out <= "01001100"; -- 0x4c
                when "1110111101" => data_out <= "01001101"; -- 0x4d
                when "1110111110" => data_out <= "01001110"; -- 0x4e
                when "1110111111" => data_out <= "01001110"; -- 0x4e
                when "1111000000" => data_out <= "01001111"; -- 0x4f
                when "1111000001" => data_out <= "01010000"; -- 0x50
                when "1111000010" => data_out <= "01010001"; -- 0x51
                when "1111000011" => data_out <= "01010001"; -- 0x51
                when "1111000100" => data_out <= "01010010"; -- 0x52
                when "1111000101" => data_out <= "01010011"; -- 0x53
                when "1111000110" => data_out <= "01010100"; -- 0x54
                when "1111000111" => data_out <= "01010100"; -- 0x54
                when "1111001000" => data_out <= "01010101"; -- 0x55
                when "1111001001" => data_out <= "01010110"; -- 0x56
                when "1111001010" => data_out <= "01010111"; -- 0x57
                when "1111001011" => data_out <= "01010111"; -- 0x57
                when "1111001100" => data_out <= "01011000"; -- 0x58
                when "1111001101" => data_out <= "01011001"; -- 0x59
                when "1111001110" => data_out <= "01011010"; -- 0x5a
                when "1111001111" => data_out <= "01011010"; -- 0x5a
                when "1111010000" => data_out <= "01011011"; -- 0x5b
                when "1111010001" => data_out <= "01011100"; -- 0x5c
                when "1111010010" => data_out <= "01011101"; -- 0x5d
                when "1111010011" => data_out <= "01011101"; -- 0x5d
                when "1111010100" => data_out <= "01011110"; -- 0x5e
                when "1111010101" => data_out <= "01011111"; -- 0x5f
                when "1111010110" => data_out <= "01100000"; -- 0x60
                when "1111010111" => data_out <= "01100000"; -- 0x60
                when "1111011000" => data_out <= "01100001"; -- 0x61
                when "1111011001" => data_out <= "01100010"; -- 0x62
                when "1111011010" => data_out <= "01100011"; -- 0x63
                when "1111011011" => data_out <= "01100011"; -- 0x63
                when "1111011100" => data_out <= "01100100"; -- 0x64
                when "1111011101" => data_out <= "01100101"; -- 0x65
                when "1111011110" => data_out <= "01100110"; -- 0x66
                when "1111011111" => data_out <= "01100111"; -- 0x67
                when "1111100000" => data_out <= "01100111"; -- 0x67
                when "1111100001" => data_out <= "01101000"; -- 0x68
                when "1111100010" => data_out <= "01101001"; -- 0x69
                when "1111100011" => data_out <= "01101010"; -- 0x6a
                when "1111100100" => data_out <= "01101010"; -- 0x6a
                when "1111100101" => data_out <= "01101011"; -- 0x6b
                when "1111100110" => data_out <= "01101100"; -- 0x6c
                when "1111100111" => data_out <= "01101101"; -- 0x6d
                when "1111101000" => data_out <= "01101101"; -- 0x6d
                when "1111101001" => data_out <= "01101110"; -- 0x6e
                when "1111101010" => data_out <= "01101111"; -- 0x6f
                when "1111101011" => data_out <= "01110000"; -- 0x70
                when "1111101100" => data_out <= "01110001"; -- 0x71
                when "1111101101" => data_out <= "01110001"; -- 0x71
                when "1111101110" => data_out <= "01110010"; -- 0x72
                when "1111101111" => data_out <= "01110011"; -- 0x73
                when "1111110000" => data_out <= "01110100"; -- 0x74
                when "1111110001" => data_out <= "01110101"; -- 0x75
                when "1111110010" => data_out <= "01110101"; -- 0x75
                when "1111110011" => data_out <= "01110110"; -- 0x76
                when "1111110100" => data_out <= "01110111"; -- 0x77
                when "1111110101" => data_out <= "01111000"; -- 0x78
                when "1111110110" => data_out <= "01111000"; -- 0x78
                when "1111110111" => data_out <= "01111001"; -- 0x79
                when "1111111000" => data_out <= "01111010"; -- 0x7a
                when "1111111001" => data_out <= "01111011"; -- 0x7b
                when "1111111010" => data_out <= "01111100"; -- 0x7c
                when "1111111011" => data_out <= "01111100"; -- 0x7c
                when "1111111100" => data_out <= "01111101"; -- 0x7d
                when "1111111101" => data_out <= "01111110"; -- 0x7e
                when "1111111110" => data_out <= "01111111"; -- 0x7f
                when "1111111111" => data_out <= "01111111"; -- 0x7f
            when others => data_out <= (others => '0');
        end case;    
    end process;
end sine_lut_arch;   